library verilog;
use verilog.vl_types.all;
entity liushuideng_0741_24_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end liushuideng_0741_24_vlg_sample_tst;
