library verilog;
use verilog.vl_types.all;
entity Dflipflopshujuliuwxwjw_vlg_vec_tst is
end Dflipflopshujuliuwxwjw_vlg_vec_tst;
