library verilog;
use verilog.vl_types.all;
entity Dflipflopxingweiwxwjw_vlg_vec_tst is
end Dflipflopxingweiwxwjw_vlg_vec_tst;
