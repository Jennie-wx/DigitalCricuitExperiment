library verilog;
use verilog.vl_types.all;
entity liushuideng_0741_24_vlg_vec_tst is
end liushuideng_0741_24_vlg_vec_tst;
