library verilog;
use verilog.vl_types.all;
entity Dlatchxingweiwxwjw_vlg_sample_tst is
    port(
        D               : in     vl_logic;
        EN              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Dlatchxingweiwxwjw_vlg_sample_tst;
