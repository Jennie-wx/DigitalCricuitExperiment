library verilog;
use verilog.vl_types.all;
entity Dlatchxingweiwxwjw_vlg_vec_tst is
end Dlatchxingweiwxwjw_vlg_vec_tst;
