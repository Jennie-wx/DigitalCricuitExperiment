library verilog;
use verilog.vl_types.all;
entity Dlatchxingweiwxwjw is
    port(
        EN              : in     vl_logic;
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end Dlatchxingweiwxwjw;
