library verilog;
use verilog.vl_types.all;
entity shiyan3_vlg_vec_tst is
end shiyan3_vlg_vec_tst;
