library verilog;
use verilog.vl_types.all;
entity Dlatchshujuliu_vlg_vec_tst is
end Dlatchshujuliu_vlg_vec_tst;
