library verilog;
use verilog.vl_types.all;
entity wxwjwjsq_vlg_vec_tst is
end wxwjwjsq_vlg_vec_tst;
