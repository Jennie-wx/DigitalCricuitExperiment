library verilog;
use verilog.vl_types.all;
entity adderwxwjw_vlg_vec_tst is
end adderwxwjw_vlg_vec_tst;
