library verilog;
use verilog.vl_types.all;
entity Dlatchshujuliu is
    port(
        EN              : in     vl_logic;
        Q               : out    vl_logic;
        D               : in     vl_logic
    );
end Dlatchshujuliu;
