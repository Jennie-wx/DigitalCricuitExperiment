library verilog;
use verilog.vl_types.all;
entity fpq_vlg_vec_tst is
end fpq_vlg_vec_tst;
