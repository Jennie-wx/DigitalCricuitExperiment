library verilog;
use verilog.vl_types.all;
entity liushuideng_0741_24 is
    port(
        \out\           : out    vl_logic_vector(7 downto 0);
        clk             : in     vl_logic
    );
end liushuideng_0741_24;
