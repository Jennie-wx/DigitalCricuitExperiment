library verilog;
use verilog.vl_types.all;
entity wxwjwlsd_vlg_vec_tst is
end wxwjwlsd_vlg_vec_tst;
